module moduleName (
    ports
);

always @(posedge clk ) begin
    
end

endmodule