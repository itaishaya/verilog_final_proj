module ALU (
    ports
);
    
endmodule